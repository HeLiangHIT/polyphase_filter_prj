library verilog;
use verilog.vl_types.all;
entity out_da_data_vlg_tst is
end out_da_data_vlg_tst;
